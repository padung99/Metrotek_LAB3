module byte_incr_tb



endmodule