import amm_pkg::*;

module byte_incr_tb



endmodule