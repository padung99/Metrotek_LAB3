import avl_st_pkg::*;

module ast_width_extender_tb;


endmodule