
module byte_inc #(
  parameter int DATA_WIDTH = 64,
  parameter int ADDR_WIDTH = 10,
  parameter int BYTE_CNT   = DATA_WIDTH/8
)(
  input                   clk_i,
  input                   srst_i,

  input  [ADDR_WIDTH-1:0] base_addr_i,
  input  [ADDR_WIDTH-1:0] length_i,
  input                   run_i,
  output                  waitrequest_o,

  output [ADDR_WIDTH-1:0] amm_rd_address_o,
  output                  amm_rd_read_o,
  input  [DATA_WIDTH-1:0] amm_rd_readdata_i,
  input                   amm_rd_readdatavalid_i,
  input                   amm_rd_waitrequest_i,

  output [ADDR_WIDTH-1:0] amm_wr_address_o,
  output                  amm_wr_write_o,
  output [DATA_WIDTH-1:0] amm_wr_writedata_o,
  output [BYTE_CNT-1:0]   amm_wr_byteenable_o,
  input                   amm_wr_waitrequest_i
);

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "ModelSim" , encrypt_agent_info = "10.5b"
`pragma protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`pragma protect key_block
m6JtfLzdUjfZ4g+RVM7b42Ls847AgBEC9h+3yJ/4Koe8OFWGkXy3nOltlqMQlNOx
avxnpqps77a6WLylR6Xid1JcPHzP64njmsul/hSd2jp+www2QHHPH7LPwpsQq25t
Slr1/hAsoqKv6/As2IphJob6sYS7w9Ty9rOXFTrIBBeFhVpePEEg4beUWgvlqgNV
ZZIzRh4aeaVec0F3TzJ3nvluyd0j8WnLzsrx3YUj4cGlWW8flKoF6xPqfblbBRQi
0yppDO/5U2lLHxfyX2OLkrOnnJorkZnCSRuiNwQKu9NVoCyECC5YPw+KK1571QVP
qebEceFx60/86LUqvW0Fvg==
`pragma protect data_method = "aes128-cbc"
`pragma protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 8048 )
`pragma protect data_block
06vHuJrLt0NpJ/6oYoORR4CK5r4l3cXy88xeN0oL0lvnqV5t4RBZHFycDkhN/57e
QyLEAMvfyloLeLkzLcbl98ILslx+o07WYyCtp73wHid/FsSRsGI0/yiuNgi1bIUn
BdYrtJ+Qy3RJ5zYZaHriXauIKBJBzEFi7cWzp029PVQth/DRMhMftyEo9y3QQr76
+49vJJTI2QqZ3F1aPyTmAokgLi45N9iUBKqFJ0aLrSFxAV1iihLwiWPtqYX3XwC9
0l7h9l5uYxQCRfdpD/EAXW8+OPkw5HudZqv/pEBhAQGzCRCDuSiXD9gIt2TDdRq3
h6ibJiqTBoVJOkIhLkJ9iJpkSEXsNlfoZ51PN4j12kLv2+aVpmHlgkQZDN2uxlSk
HIIhucQdaTSWw5k/tCYx3a0n9sB/1qpec0imtyDb+4I4N2daqG+yoGuXqyjqrONY
HlkcBUymebFfxx5/qhQWKF9jSUGqtMXvPrdWIzRaofvVktJ4wwQglh5ok/S57NM/
G4imdJmH2Zdpk4ZTsTfMIgGRNoW4gmhIZn4OyB7O+dPD7w0B0DnrIWkVxKNLxIXx
nwnmUwmXcC/ULds4rhtQoczQzmPD9GBEl2L8l9ehoQcI6DaQCre1rdwGSzwOi6DN
BErgqTXMoqBLi//oYx/aHre4Y3j4wd5WWhaH8oragE/y7O3v/ngnEK7aKrz0Sp7C
bcfMWsca/h8iY7PomjVNTyOoGChHBiyFU2/5SL/L70Y+swlXMm9cKTE/OhkfNPPx
kt/0GWx1PIIUrbbJRLvd18O9xsDFXoRISPzfabSq1XhO93nbA/w3davAu+OH/A1Q
BQ72MPLuzCN+xEzSa4UHGwrMv/XYQU4Tq3Incig9D0d4j6oIg91qngJxapO0bmKn
r3XGCpXLDDFNbguRDCig3m6zW58eOFuxzQubsdZ3gHEC0yFg6ffOz6mJsyg22KSW
5x9KcjgtvZFpGFKceSrDJZwCJjCiJMEZ4htahADmM0ZsRajogoJXw/YOR94RDM55
OCQwSx3+0YpH42D9bnvY317I5LnV3UBOQf0I1lthnpy5tGmp11rcm+XpUKtuvSJP
7KZwo+zV/8fn6b9UmOpC9TNWkOABsB/bbkJPCiGQ3gx46D0Hdk7tP2gzFyCcIWMV
SSpJTdKQhSQ9Zu8kSI9PSNFUwSZUE6Y1zVu6WTirdGyOX2QwlzM2FOO60kfH1N4u
BwFk9t5XODIBDvrDFN4dGC0edbvRUiwc/YSp/e9o2XT8cUAWNjAfUS+kCrgOrSZJ
Ff+b1maaU/MeAzh4e4xMiSeil3/hp50Xn5Ffpg4IgoYW0d0czs11y7PB1WXl2z3K
Wf/MSvM/AHpL5oWQ1MzruhSINzGJ6E/fPyAe6Oinz7RwMU+0lYeTOMKz3IO1UvCw
Ak8hlHkNiCEr8rMmZxvfwWd2WA6cNJEERYESab/3dUHqi+vjxqaqKjsvvGin+gMU
tqNmV9dO2r3tpn3m0Bi5t58vXTB1DPGtqgnxn2QkdyAqzsM2flY4krF+ZPJxuDN4
0fM+1mf/pvoYB5tuDtovN364FSsCqVK7fh/zX7o9tSfyRblCd3wtaeoiaZ3vrqQO
Dztv+P52fJ7G2LYmW2K35b/dSHUHg09miL8Imy8RX4E57NAS/VMHAJ4EfKUojooS
BwUE3IVHTMkKzwS/OfrlAu9zlHXF3SVmc/FBkagsptwiDpF4XQciSMR24g1wodAs
pkfBPIzml8BtdSnm7O0tlNt+4U5V5fl6XizmtiZxjg1CgcFLeI3DuPtIufS0rf1u
zfYhNArPpBNpehgAbZAMVqVKL5jtlmp5blx3EGgGOu0SFCfRZ69Z8R/gF9NGiCbm
h8XhRvrv9ourqbyUg7aOXqN/DxDKTnEmPlRoY6Pf+EEGaCwCehJubGpJFoRzEjMs
g/TIfJH1jAhm330etqvlANQx2z3JW+9dyLlG9PXQm+Ikcb0bznu7xoDr8tMJWKd+
LnIkNGOrWBcWFxFTq7kjbaAtdaj1zyqCHwcaC6H0a9Ui2EH9OrfF0YCMwDXd8AAk
XjK64QBMpHcOJ8eGskM0BRJIsbQq9gTuuPzmWunKX0KyaURyjRJyhdEKVKul+I/i
YgSsQQghsWs1Ab62QnLphvtVMN97h3lnlvRtmCTpXdfW7497GwYScKVWm4ISWsDe
zB9TSyrxk3ogkp293FQGwvbGxK5YXol62hwps2u8TH1zFM9qG08hyRScz9O4Tws5
iRBLP8kY+07EvFAvqCMa7GKsJmI/I7oNvM/bUvAKD/1edijBoJU3c9GZrgYr4MjP
HIN85mPc/LRq9fY8VwENPI+WpijldkdL2OxffQiwpOAzST+4/36lkVJF47eovTeZ
wj0QbtIPn95HdvxcELnr5qVYJmIgV4tRXEdi/KhzepO357WL43/ycau+BWl3Czkd
bK+0l0f5AzJGmgKujxXFdX41Fm2gVkaJ73UVdXuMqTU12hvweSuZxf1wODi0QFz3
bbvsE6UZ0GP5vk8eTf9rA74urar/xYB3Ka2oKukt5ru5eD1EOORtzMt7Re+WA2A7
D9eXlnXhmOKebwIO8LLXtyYgQoAHG2WCl0bq0L8VRa85xc7bVeWzLHLmgZ9cnO40
RWxWvZHSGRCKUshviudo3y5NHeaQisTNkg5VUYkbI5KgGzfB0168DY1emUdJMsL3
gy3F/FngSvZCSiLJ81/j6nomCTPTkbAmSnG8B9ExBJTnIrflpxateDo7DklKP/tz
NyGAcYyBfEtMKGKC/MlibkP7I29GeiEmaLwvPazyX8eHASDJvuxmS3kWIOzd0aEo
/rd6WQ1MEBriXEjbB9YxXehA1v5GJBsrhxNl/2G2kOopYGj8RxTpMDAhb99GYQdd
Ar35XEqavEYU4t4KBXObvaFZbQnGFIzvGcIFIF32p9oqsK/lyK4aadi4Oano4y3y
vVpTBRsAAzEH5yq39KFCnYwiqXiLW60wahmBch3ygsMys6i1aefEmofI4eQfzX2n
NL1JuM/FE7soKTpYy9kKKfS+guIiCSpwdbSYZ1Fxy5ui/n8jc97y6TlCcOgdMKPR
kIWVboglT50vYke8YbgYwA2DDWad8UjStef0U9BJxb+/VyXpjDf6k49ZNz/Aeuwk
9tf6PqFOydSoQuykqvYU1DklE+ye54RoMEijuuI6zHBnhkmCrsgZ6Q+XLy2o8mrz
twZ6PJN4A4QH2P6I/ky/9w9sW6rq1Nd7S1BNTIfh2tPBL9mYfucWG0EBxkTRkOau
ISkrLoGmtcHEOBNi7fVYhezNt+F45ior3MEE+iZ/94LfvIwX3iZIbTxgN7PSldEV
WnOu4zSSzFqLqEEYW4aeLQbX1BT6RtVQkFDhKhQwWeqzmUdiz3YZQHOGB9FF9eo+
bR3mL8MMRnqxFxZ91jF1rOn25IEiClUNwnJTLDjygXu2oWjpYxNVapSvgwoZroJG
1w2jKm0XXEWNw5tB0HW22n1NAhVEC5ZmIjBgGhHMR01DIVj3J5hq5er8lS/DPpCh
39vZoTir5Eka1Al61tAoEm4w0FS4WQ4bQxRpZjWQZk3dGj42DdTmE3bGZCoEkcnn
INiKt8MqP/AKGoCDCWgX9UqGzNgDEeqwVKYfo7rIlKhWQnEb0yUgl6pWMsm1BO2W
U0oC8xzKBCS1+ewBZaF2NiSWLCCslKzXjIImSQBo0+7lAFG5Z0M2yyAnWtpLXnql
7boDRcGjy10Mf3AQnUtgio4LgHDhCUvXRut/OGKV2X7hLUf2w4NhXVNCNbU1RvoX
o7fyz2p+IGffM4mk2YOjksO7AScTH3Pchwtk6fhnO4+5qmjvxvu8wkNtXMelh0MR
IqalJ8LlaNNAtQ068QpAASrvGCez6dRWGOc5OOaLoY1vnmngz5YuOhhLgn5uCmNF
rIgjqQvrm+lXO7VUbe3gJoNewfoeDjgitHsLvw2EUWzXbofs6ZrsestoqZ2WkkIV
niQWs/PRt23w+SoamXefJ8YtAbk81kyICE02SkUvwv3Dr0bIPNTdRVy+9UIivZ6G
dDVEowGuqeXpj8C7pLQ/lpuJgxJKVZBcCNEGTkVN/3Rtpzmp8pLA//oNYmGyWbEA
IljfTkJCojqpi9VuYsRbRqstjxHtxB62CrSivWfToRgO/jE3MI9s+JVVUyMyZstY
yIMoxnRgESiZ2Nn5DXQ8470hctNeNGmrlV8serPMzHXIjol+hvdu9o+Zk7/wmvMO
DSB4SIc/24vKgbsWpDSHsqg57SAgiypvcZVXVtq/mP1wJSL6aJ44V3NbcbgFI8+J
MtX8l6jCuxx6utqhw/UvLuSHfsCPF5H1s2BZ1cZ8lBzBwNJAzW9W4hCB80cyyHw2
8qUdgI5JWeyuVDTf4HJ/TBLjMsPm0ffY6lvBzD7rluek+fKjfX3wBeIRATtND7Zt
U0eHPlX9fv/sgAgtnrmmmwsj0VuiN+Gt12YdNOyzgYOWTkrMeFNZuKYeJumRuIgi
Im+2t3h8/lf59qDHD5PKgZUVxG7X47knXs713/O987pp9LCQowpiSW6SCrad6zem
Q3acE/VN99x1WsuIzPZweTcUsB7BOjHBb1XsbcPP4occ4/9sYv06mVXe4Vg2Phpm
Tb+H24u5a96MGx1uc7gWxScppZ1YmxEFqDLJgWjOMjC5+L2SUjr6/n+xqdVrryoP
mTPtvIQLwsc2J1CNez86srWv1hhs6xfBvCIVKDa2sTCB3XkI5NK2g3Lx5Sy+D4q0
hW4Z9yx1cQpnkYOJ+qVcr91BtJXiW2SVgeA4RhmeGF1eo8sA6QhsPS2/t0gIzyet
rkspHFoncRpy2cD660jn91pLsFzSNUh7Enzf19V42/QLoU/IDWTxT8l9eMtKVD2t
UO541OPYq/nDzJBI05oJkYDlCK3OKc8WNb4wFD/iTryRZNEfSC22UO90YevVoR3v
Pq7CIblYQtVArvC3tiePqZf7JtGBvmhhEX8GXH2XV/5iXeP45WbhyMwMx2gYLfOP
+v7cv6OH2A+CzF8V0BiNY9m6l1bew4QZaK76wvAK2jLydwROKi9G+2ahwEMlpZqJ
D36+3D4Zii1nlHBSkZuH+OruaP8JZHLM6vWZfLWbwI6jmXDu4Rn85DF1gNK2Jtlr
qSJnxu6DUm07hlzzEIkuNOVBgSioCiW4T11IqCXAA4ASb0dzVl0nZzoHsjB49XzP
NMSQMw6eOcT5hqhxYGfWtjfY9qA6YbEnzCV3OLtdpMX1wjX34loXidtoNgPngT02
WkV9qJwTrbqBqrrzEUV8MRgkc2VhEc12UUwnzZODHcMCDRPQQVj22CCB1QS6OUrv
3NkL/uxTmAM0QqVfuS26hzHrC+vmBZOPECvLNNQEl7npOEWtWm6xt8epvvtOlfNM
nfC+d1wyUXKaMAAjbzWAJ+bS/QoSivm57r0Niyh9Jd14Kwjvy2nCgOwleDdt3RxO
0ZxWyOXULnY4TD0zZDcm/gvIElRvdgTBv4+vNWcv27nx3GDYzAMU0b5r8aD9MMrc
q1OO5HaXOaBIQ9z6ctXDBlIAoqLRO1tDrzLCy1rSlHyNAmQ4UDbHomgbT0oPCgm8
SPaOxhMOaSwP525ci4+WzujIEIH7FDGY0dlJhG6TKjuf6AXRohFppMCu/zg03jdO
1pAd6mvE62H9mohEnup8PR9uUerqUcVCLjlboEPn4WfPLG2vHvnBwtll55+L0EaD
9hILLeTm8/d3U55Uw7pngMti90DMuCofL2wi6iVsWlbtafI6Mv6Pr1GWdDUIoel+
ogfjphtFynYu3vp9CNCUfJr5LE6RKY3ByEy+TKYXG5QkwgXDCxKCkLJIYHk/7XmZ
ypTp6CRDGHCFevXEFDCZIN0/YA8Gu9lAcoIcPXP7b6jZbW3dbKUZDp5pD71V0vfy
X+7VGWKVxuf/h8NXfEOGWtuaN9ZIenPIm6rV10mQjXDV/5YhlvV0CYis/h7J4k+z
8s6UFOrA+Pc9iiPFLQvCN8pqhzXeHNqYq631eSaUxb+NYIireBzpjXQzoQjwSQbS
z7vK+9b4P+8dGGfhX6yrSLkO46tuAwYSsFIGSJmZNoUqakfPDm46f9hXzyisUljz
apBhEDBXHs8i8cnKn42rwgP0nyQWKG7+JIiYghujxjWwQpt8hqbB4Q0KJCF9OiUH
eJeKYPWuvuZ6mbT7oId/h7/bllZ5jDUb7vIADazoNTJQ1D9+VWmJf0Cwb7+GsIhz
HABniGkBU2ShkcN4BuSmj0rm+geFQ2PFHT4OPIT9+0A9DlxFRyotQgeEKY5HHN0R
UimgwbagScTiehZJB+uqOnbDpUYx8d/oEfrp32rKmLRDssr62J7wQIgryDob65ep
gOx/IFiYxgc+SJmXEQ4cioQTbvQeoSAZTSBnL8YQHoJlLBASupEIoVnbd3cUpVJw
+hr2roi5DKzGM/te5Lyu8pPMy+Vfkel/uq6vHp9h3+6gh45/5Jzx/u33k9QN/eD0
qnlDVBQciSJ1XH/b2HzVPOKWfogkdAqsQl5GanDfaDDQS1fU0yG4mJeGzGtuiXlv
O/V+v+5cNRl1w8qDu43FAGoPRNKjklG/ScXiRlBpdt3SdrHRP4NEvvq6jH6x1tPi
jHyD/Hz76yibq0cjcrhkDxz1IvB3lHJNb75skhNUdGQeJ8LE4uR+xivABHNGzhQf
JIlQBSaiRopNHm0QuRZpVSJIALyD2VtTd2Zx3sSa+8PhfSYfHJtuNjML0pBufQDQ
07Xl1TbBuhdYnKWX3Rp73U0pJhInpUNJPtr1nOH+m0QKdw/NwMnL+QTbC4D1nETC
Wcu/VCUTXY3A53BMN0JC5csKgNTUe0Jxh6nRUxXudB5tfqxr6xBVbRKJe7EMbnmT
DddV89KyEiSnMJSsl8drkB3eTwm+IIfmPnT9hJK6SXf2QFoZN9J0TY4hmlcjLE0A
6DVBV9KDZhVrH0tKNubHK7P6fYmLszqCJ6m0NjXh34TTgXcJPFpmRw/bJw3NWrrw
LH4Up+/+VZYqDYLbWG2m8KLB8iAM9GJ5AWFEJlIxp7Ji6blcrnOs3o25ufQm2LUn
F0dg41lzV2dxzmAHWKe2kXMgYwbfv3WNIK0ODnTvf0HkLQzJtq5SqFzfe+LA9pJp
cAIEXh3BUUM4g2JNbYFnd4kwUVAvSIrtnnAh3VljEDIkSUe9mPRNsc+O6DGYzVxk
lbjI/CufTkQ8wMvWBfjLI8jFoxSf++c+TjGEGRMnhRDSXWUyqjG6EtirA5NF2bKO
JhmqSvAbIeH1n+KEbOLPPmHjGwFzDvY5V5u2VudcyIDxrUjdFcDd8cdKC92zn3sy
x4ZPsZpy6Nax8jBXbmNJS1QQzQzKZy1RXTDmtZWDae21w7g/0VjwyzliUP0+OMmD
sRI2KfIqXO6tSe48f0vSQ+1djV0/N2TC3U0+aOL24lwKJ8ettIlZMv0d9RMZkJ+C
W7aU7gMozi/Wyq0Z71hvdDLDJxFa9XUSuZmQC98SE9HJDNv4FfW6iNSL/s/RR34s
efnV3iBOvKE/fm7hizH4E2tAjFSX5a01fImxVXcLJOk2Cnpu9ayU8mxPvbDgYGBK
2lxxv2n/gdkEMFNXgUrsCc6ADkWfODaCxF3aKt5bJxf6ig/9Tm3KK7NkV4mS3ho+
GLgQgZzxhp872OeAnCuSXVMWI5zaBr0PoY4usfT3iKOCg+e1cvHYD1R4XJxWg3hw
8n+tdcsi9pcIW5pbikIofGly1F+sdnri2C/HLH36R7VOtx6Ml+fdmThGeerb+rwM
Bn4L/13pVv6yDoxrN8rtUovWfZGiYB+1zalrkkd4YxfUGUA/fWwrx2uejAzMs7iG
A9QLWU9h06haN6UDqcWNpmO6od5yBsuucz0h2Al7AmB8Lx0WDc4Jg+eK0fdvBop2
91J/bro5tHUav1uHa0YtExQSYn98KfgcEn2OKPAqtII1iQTi5ms5Qv3UgL2UQHa2
wTXbRuixYZZ4/sl50C81HpxteiUvlFLVTsCzyr6yvYDjUCbrO74GGS4BXYl4ZtxU
EoHcvF8r38FGIrtmbLxDag0jrzCHHJPiQ117x/chYN8lLWRWM6LfkajcKHuFssOZ
diTxs7X7qf8A3tecrVTeirCktL0pkT8fTETGK4ogk8yedlCLZrMyptASK3H7O+Ws
Jp6q6TAv9zE20NfmDzdain+GA+aoU7PvGxV86TXI+6w2FLeICj7CCWm6z2hTNp7p
73rHVYzj8SFIeM4rWGb/FqNzh5RlS9ygNoh0CvEnl7fimfa+OL+BwZ7eTcSbJI6V
2JUCmndwSwlDJDF100yqSGQ1x1axHC2PA9nNUYAkeUeE/51AJqT/r8ukHNM42Dq9
OalRQ+gWUZ6GklZosQeezHbPJkDiHEd4icpRdAhWicDVd7RoYencKAbUYVbru1Wc
T7/sFRbkG0SOEvxuYRJLlHsbizqsdwhjOrk/KaTgsTd58n0O/tCtUzEBSbBJenJ2
VOCCYr3HXtRcEtwkze8Wola5p6vXddergR6/LughaurEg2hF5cSflyfSZj2Ww6Zt
0tFkQ+0mFlu6q6TbqSXU4HbKXj6FKu7pFpSN+y2UnQtVDNCkCA9fTRkwkqXl82Mr
gDdRrWMnyomyGEaYAhPALXFa7cEzfNUytcN9e7wWTSbV59Y+baNIToLH9Mjmqmkv
H6ImZbMzccV/sxnx5kbeJzsMLIfLYu4GXsrGHLeUhoGtVaPc8I11KNyRIUsaEBol
Qm7NTJho64oAnE1jMdq11d9omX43z8snGfgaWGU5M5fCPam9pt/Tv63uYwT2ckBZ
tCrGpe2qcoTa4Uf5gY1r9GzHhAToeg5VOTbC86jxNUJlP2EyIm7VP0zDJxeMaHR8
jTwBGVLccHRlRTYQ+WSQIlwt+YwmDEsuDVN6FPLktesMGNpwx+NW/UDacLyUUUi3
wfh0fE3/hAtMpTQANrSM00uV6C2hb4FYiytSJjfFwDO6Q1T19wV7lP9rWxKgjbs5
VEfTENSGIYupJtTMBTD3nq/ZvYMbm94iD3r8plHs0xacSg+TvCR71I8Rhh0onQXn
RGs0dH9MZrJgEWjST/rBFpT6gIFMDs4PbYlvf3mvFwzcMdspWTo02xOqVhAoD/Gt
4w7lYNBcH/u5NlRWLDYT3jIRBxlcLmVX7Vn5apDqV0Z1jMGXRnIYyvFA0ruahrYS
dbs5JDa1lxuwEh5gljFA+SELyfIVTFScJhERfkqfqGzHIs9lMtZK14IFFQ972qM0
5aOPr00UbLNw2W8OYL2NMgExYTUlO+6ZZ+O+lh3MxfcQOr/FwXQb6YNceDsMzecA
0G+4S0/ua8dWTfnS1fFBSXUVGlIDVEIPOIwVvHqPpTMenOwGXuy90fg3ifC2vNMz
QZFEcw3JVGv3rYgDlwf189CTm8i9H9oAfH91wERIiZIGGi0LyVQjLOyu3kKVyXBk
ipgtpTh4NlwfsFqcGn6WadtLZ6o1xP4cppueFkqClmugvfbbn0SmzbFKecy+spYo
GmwlfYN/G3rTHg8sRptXEzSgKQz8cKv622SCoivs4q/fJ5v92QfFBd2stf0Nyk4J
VnTSZYt6YadZby5s1IrkOcAh2SmN0HH4OCKY+KI8xtv4Oq0dj1B0Jrszm0/El6PR
sSAcAZp8SnkqVhtTEI44Wo7JIaZpB044aGS4Z6CBrZSb7kFg8/hDujD1skyHaKLt
nUM+lmLw+rVB5C9KXrn+aPxNv6DP4FUADAtIHpgRHIXaIJwmrelVG9fd++kfYuX/
IGGG+eVdRe1zE+x87t9lFu5dl51DNrGzpO5XX++kUIKzmPYjozNDXLSQo4AeEX1x
jQvwnYJT3Estjl2Shn/bv1thUExPX+cn6cAm2gu9ZZgr0Cs4YklgUR6erQa3ZIXT
/NY4Q2kW71ZzsMq72clKJ6+O1m+7wsqypzlaDjq6WaPDok+q5/7zohLwAcBKDxh+
127LJJbmNbTzEwM5YVENA7HUr08KEQ2ip4qWSWju0E3XBgfVfLU8BEidS90SF+Ti
qo1w7wxoJP4QwYIUKtrMusI7aGb1Eb14+d0E2NXSvI9T8MCMxnq8UiAa5dEEDwGQ
QQKFqEL2oKZtbwOutXZBVFrlUHAIene+FCk0lnrD0PTria3Q9msRuAgbrBetCxho
dKNRrXP42Z8k6Uvs0DnUibYs5UzUJXyUDnG1JibVw2VAHgq9OwpIVXm5um+y+2h7
2JcUjqn5fHKyjMsNhhCnCAd4ebz9iI5cTiZx6cTi7PQxArvcPd71ajL+k347Sgni
F2C2x0wwec6ZnbIGj8WoZC0/FaEiMUcz2j36/amEjkcyTRjDwbZVFEypiplEQ31I
Fka7WkU/t5JoJhwDV/9ngLDyY08JZCFS6DrO5zmqZ2W7DsDHTBrqlI6ScNFTGF3N
2TeqIFcYpFlcileYyBgWR8MrbTJUtKL31GuMmvbtJQjgt1C1Xd8RAiNqS6LQtFeI
s/wXaBIhGVnNRe7L8Gp3TJlGvoyq2qsdxmUSRkqjeuuZXwSPTVpZ+g7cZ637r66q
bBXwBCKjZLV2njGTSOUHekjnTiQs4q4DAV2cqedqeViJV65efvrHA8YtHctl63CO
T3TJyLbPNKN9b8XSseVebaf9e9pdgBzzdnSji89bn7ZYqpZYAaF2DnjipGjEx8S9
dIqpjGBzdmIfMnyGDuWo7t5IbsUAi9MGC51df4/rgOOOfCFeSK6OuOph0eH6GLeF
jTUAaQ8d25myYYniRymhKDDpdJOCTXANymFRMLwSU48=
`pragma protect end_protected
