module ast_dmx_tb;



endmodule